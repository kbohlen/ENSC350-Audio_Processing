library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all; 

package BandPass_FIR_package is
  constant SIZE : positive := 16;
  constant TAPS : positive := 57;
  type coefficients is array (0 to taps-1) of integer;
  constant C : coefficients := (-904,
  1503,
  -5130,
  10246,
  -19998,
  38213,
  -63275,
  106688,
  -165043,
  251083,
  -365383,
  518408,
  -711779,
  954562,
  -1248331,
  1591847,
  -1993118,
  2434750,
  -2922821,
  3437740,
  -3970909,
  4499114,
  -5022604,
  5487076,
  -5921931,
  6264614,
  -6520104,
  6699513,
  -6727994,
  6699513,
  -6520104,
  6264614,
  -5921931,
  5487076,
  -5022604,
  4499114,
  -3970909,
  3437740,
  -2922821,
  2434750,
  -1993118,
  1591847,
  -1248331,
  954562,
  -711779,
  518408,
  -365383,
  251083,
  -165043,
  106688,
  -63275,
  38213,
  -19998,
  10246,
  -5130,
  1503,
  -904 );
end package;