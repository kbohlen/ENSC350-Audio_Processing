library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all; 

package LowPass_FIR_package is
  constant SIZE : positive := 16;
  constant TAPS : positive := 61;
  type coefficients is array (0 to taps-1) of integer;
  constant C : coefficients := ( -43,
  38,
  -169,
  174,
  -470,
  524,
  -1073,
  1257,
  -2136,
  2588,
  -3829,
  4749,
  -6302,
  7938,
  -9645,
  12264,
  -13847,
  17683,
  -18764,
  23963,
  -24115,
  30677,
  -29491,
  37236,
  -34408,
  42969,
  -38368,
  47228,
  -40940,
  49499,
  -41832,
  49499,
  -40940,
  47228,
  -38368,
  42969,
  -34408,
  37236,
  -29491,
  30677,
  -24115,
  23963,
  -18764,
  17683,
  -13847,
  12264,
  -9645,
  7938,
  -6302,
  4749,
  -3829,
  2588,
  -2136,
  1257,
  -1073,
  524,
  -470,
  174,
  -169,
  38,
  -43);
end package;